`timescale 1 ns / 100 ps

module tb();

reg clock = 0;
reg [9:0]SW;
reg [1:0]KEY;

wire [9:0]LEDR;
wire [7:0]HEX5;
wire [7:0]HEX4;
wire [7:0]HEX3;
wire [7:0]HEX2;
wire [7:0]HEX1;
wire [7:0]HEX0;

top DUT (
        .ADC_CLK_10(clock),
        .SW(SW[9:0]),
        .KEY(KEY[1:0]),
        .LEDR(LEDR[9:0]),
        .HEX5(HEX5[7:0]),
        .HEX4(HEX4[7:0]),
        .HEX3(HEX3[7:0]),
        .HEX2(HEX2[7:0]),
        .HEX1(HEX1[7:0]),
        .HEX0(HEX0[7:0])
        );

always
    begin 
        $dumpfile("project3_tb.vcd");
	    $dumpvars;
        #20 KEY[0] = 0;
            KEY[1] = 1;
            SW[9:0] = 0;
        #20 KEY[0] = 1; 
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
            SW[1] = 1;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
            KEY[1] = 0;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
            SW[2] = 1;
            KEY[1] = 1;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
            KEY[1] = 0;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
            SW[1] = 0;
            KEY[1] = 1;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
            SW[0] = 1;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
            SW[1] = 1;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
            SW[1] = 0;
            SW[2] = 0;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
            SW[0] = 0;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #10 clock = ~ clock;
        #20 $finish;
    end
  
initial
  begin
    $monitor($time, "clock = %b, SW = %b, KEY1 = %b, KEY0 = %b, LEDR = %b, HEX5 = %b, HEX4 = %b, HEX3 = %b, HEX2 = %b, HEX1 = %b, HEX0 = %b",
	         clock, SW[2:0], KEY[1], KEY[0], LEDR, HEX5, HEX4, HEX3, HEX2, HEX1, HEX0);
  end

endmodule